// =======================================
// You need to finish this module
// =======================================

module si_alu #(
    parameter PC_START  = 32'h8000_0000, 
    parameter INST_DW   = 32,
    parameter INST_AW   = 32,
    parameter REG_DW    = 32,
    parameter ALUOP_DW  = 5
)(
    input                   clk,
    input                   rst,
    
    // arithmetic
    input   [ALUOP_DW-1:0]  alu_opcode_i,
    input   [REG_DW-1:0]    operand_1_i,
    input   [REG_DW-1:0]    operand_2_i,
    output  reg[REG_DW-1:0]    alu_result_o,
    // branch
    input   [INST_AW-1:0]   current_pc_i,
    input                   branch_en_i,
    input   [INST_AW-1:0]   branch_offset_i,
    input                   jump_en_i,
    input   [INST_AW-1:0]   jump_offset_i,
    output  reg            control_en_o,
    output  reg[INST_AW-1:0]   control_pc_o
);

localparam ALU_OP_NOP   = 5'd0 ;
localparam ALU_OP_ADD   = 5'd1 ;
localparam ALU_OP_MUL   = 5'd2 ;
localparam ALU_OP_BNE   = 5'd3 ;
localparam ALU_OP_JAL   = 5'd4 ;
localparam ALU_OP_LUI   = 5'd5 ;
localparam ALU_OP_AUIPC = 5'd6 ;
localparam ALU_OP_AND   = 5'd7 ;
localparam ALU_OP_SLL   = 5'd8 ;
localparam ALU_OP_SLT   = 5'd9 ;
localparam ALU_OP_BLT   = 5'd10 ;


always@(*)begin
    case (alu_opcode_i)
        ALU_OP_NOP: begin
            alu_result_o = 32'h0;
            control_en_o = 1'b0;
            control_pc_o = current_pc_i;
        end
        ALU_OP_ADD: begin
            alu_result_o = operand_1_i + operand_2_i;
            control_en_o = 1'b0;
            control_pc_o = current_pc_i;
        end
        ALU_OP_MUL: begin
            alu_result_o = operand_1_i * operand_2_i;
            control_en_o = 1'b0;
            control_pc_o = current_pc_i;
        end
        ALU_OP_BNE: begin
            alu_result_o = 32'h0;
            control_en_o = branch_en_i && (operand_1_i != operand_2_i);
            control_pc_o = current_pc_i + branch_offset_i;
        end
        ALU_OP_JAL: begin
            alu_result_o = current_pc_i + 4;
            control_en_o = 1'b1;
            control_pc_o = current_pc_i + jump_offset_i;
        end
        ALU_OP_LUI: begin
            alu_result_o = operand_2_i;
            control_en_o = 1'b0;
            control_pc_o = current_pc_i;
        end
        ALU_OP_AUIPC: begin
            alu_result_o = current_pc_i + operand_2_i;
            control_en_o = 1'b0;
            control_pc_o = current_pc_i;
        end
        ALU_OP_AND: begin
            alu_result_o = operand_1_i & operand_2_i;
            control_en_o = 1'b0;
            control_pc_o = current_pc_i;
        end
        ALU_OP_SLL: begin
            alu_result_o = operand_1_i << operand_2_i;
            control_en_o = 1'b0;
            control_pc_o = current_pc_i;
        end
        ALU_OP_SLT: begin
            alu_result_o = (operand_1_i < operand_2_i) ? 32'h1 : 32'h0;
            control_en_o = 1'b0;
            control_pc_o = current_pc_i;
        end
        ALU_OP_BLT: begin
            alu_result_o = 32'h0;
            control_en_o = branch_en_i && (operand_1_i < operand_2_i);
            control_pc_o = current_pc_i + branch_offset_i;
        end
        default: begin
            alu_result_o = 32'h0;
            control_en_o = 1'b0;
            control_pc_o = current_pc_i;
        end
    endcase
end

endmodule 
